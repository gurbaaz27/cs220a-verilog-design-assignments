module process(valid);

    always @( posedge clk)
    begin
        
        case (valid)
            3'b000 : begin
               
            end
            3'b001 : begin
                
            end
            3'b010 : begin
                
            end
            3'b011 : begin
                
            end
            3'b100 : begin
                
            end
            3'b101 : begin
                
            end
            3'b110 : begin
                
            end
            3'b111 : begin
                
            end
        endcase
    end
endmodule