module process(clk, memory, state );

    input [31:0] memory;
    input clk;

    input state;

    always @(posedge clk) begin
        case (state) 
            0:
            1:
            2:
            3:
            4:
            5:
        endcase
    end

endmodule